--register to signal map table from Document Version v1.5.3
 SwRegister_sw_HW_ID  <= swreg0(31 downto 16);
 SwRegister_sw_HW_Version  <= swreg0(15 downto 0);
 SwRegister_sw_HW_BuildDate  <= swreg1(31 downto 0);
 SwRegister_sw_ext_abn_intr_src  <= swreg2(31 downto 16);
 SwRegister_sw_ext_norm_intr_src  <= swreg2(15 downto 0);
 SwRegister_sw_exe_cmdbuf_count  <= swreg3(31 downto 0);
 SwRegister_sw_cmd_exe  <= swreg4(31 downto 0);
 SwRegister_sw_cmd_exe_msb  <= swreg5(31 downto 0);
 SwRegister_sw_axi_TotalARLen  <= swreg6(31 downto 0);
 SwRegister_sw_axi_TotalR  <= swreg7(31 downto 0);
 SwRegister_sw_axi_TotalAR  <= swreg8(31 downto 0);
 SwRegister_sw_axi_TotalRLast  <= swreg9(31 downto 0);
 SwRegister_sw_axi_TotalAWLen  <= swreg10(31 downto 0);
 SwRegister_sw_axi_TotalW  <= swreg11(31 downto 0);
 SwRegister_sw_axi_TotalAW  <= swreg12(31 downto 0);
 SwRegister_sw_axi_TotalWLast  <= swreg13(31 downto 0);
 SwRegister_sw_axi_TotalB  <= swreg14(31 downto 0);
 SwRegister_sw_axi_ARVALID  <= swreg15(31);
 SwRegister_sw_axi_ARREADY  <= swreg15(30);
 SwRegister_sw_axi_RVALID  <= swreg15(29);
 SwRegister_sw_axi_RREADY  <= swreg15(28);
 SwRegister_sw_axi_AWVALID  <= swreg15(27);
 SwRegister_sw_axi_AWREADY  <= swreg15(26);
 SwRegister_sw_axi_WVALID  <= swreg15(25);
 SwRegister_sw_axi_WREADY  <= swreg15(24);
 SwRegister_sw_axi_BVALID  <= swreg15(23);
 SwRegister_sw_axi_BREADY  <= swreg15(22);
 SwRegister_sw_HW_ApbArbiter  <= swreg15(10);
 SwRegister_sw_HW_InitMode  <= swreg15(9);
 SwRegister_sw_core_state  <= swreg15(8 downto 4);
 SwRegister_sw_init_mode  <= swreg15(3);
 SwRegister_sw_work_state  <= swreg15(2 downto 0);
 SwRegister_sw_arb_check_en  <= swreg16(8);
 SwRegister_sw_init_enable  <= swreg16(7);
 SwRegister_sw_axi_clk_gate_disable  <= swreg16(6);
 SwRegister_sw_master_out_clk_gate_disable  <= swreg16(5);
 SwRegister_sw_core_clk_gate_disable  <= swreg16(4);
 SwRegister_sw_abort_mode  <= swreg16(3);
 SwRegister_sw_reset_core  <= swreg16(2);
 SwRegister_sw_reset_all  <= swreg16(1);
 SwRegister_sw_start_trigger  <= swreg16(0);
 SwRegister_sw_irq_arbrst  <= swreg17(7);
 SwRegister_sw_irq_jmp  <= swreg17(6);
 SwRegister_sw_irq_arberr  <= swreg17(5);
 SwRegister_sw_irq_abort  <= swreg17(4);
 SwRegister_sw_irq_cmderr  <= swreg17(3);
 SwRegister_sw_irq_timeout  <= swreg17(2);
 SwRegister_sw_irq_buserr  <= swreg17(1);
 SwRegister_sw_irq_endcmd  <= swreg17(0);
 SwRegister_sw_irq_arbrst_en  <= swreg18(7);
 SwRegister_sw_irq_jmp_en  <= swreg18(6);
 SwRegister_sw_irq_arberr_en  <= swreg18(5);
 SwRegister_sw_irq_abort_en  <= swreg18(4);
 SwRegister_sw_irq_cmderr_en  <= swreg18(3);
 SwRegister_sw_irq_timeout_en  <= swreg18(2);
 SwRegister_sw_irq_buserr_en  <= swreg18(1);
 SwRegister_sw_irq_endcmd_en  <= swreg18(0);
 SwRegister_sw_timeout_enable  <= swreg19(31);
 SwRegister_sw_timeout_cycles  <= swreg19(30 downto 0);
 SwRegister_sw_cmdbuf_exe_addr  <= swreg20(31 downto 0);
 SwRegister_sw_cmdbuf_exe_addr_msb  <= swreg21(31 downto 0);
 SwRegister_sw_cmdbuf_exe_length  <= swreg22(15 downto 0);
 SwRegister_sw_cmd_swap  <= swreg23(31 downto 28);
 SwRegister_sw_data_swap  <= swreg23(27 downto 24);
 SwRegister_sw_max_burst_len  <= swreg23(23 downto 16);
 SwRegister_sw_axi_id_rd  <= swreg23(15 downto 8);
 SwRegister_sw_axi_id_wr  <= swreg23(7 downto 0);
 SwRegister_sw_rdy_cmdbuf_count  <= swreg24(31 downto 0);
 SwRegister_sw_ext_abn_intr_gate  <= swreg25(31 downto 16);
 SwRegister_sw_ext_norm_intr_gate  <= swreg25(15 downto 0);
 SwRegister_sw_cmdbuf_exe_id  <= swreg26(31 downto 0);
 SwRegister_sw_sram_timing_ctrl  <= swreg27(31 downto 0);
 SwRegister_sw_arb_weight  <= swreg28(20 downto 16);
 SwRegister_sw_arb_bw_overflow  <= swreg28(10);
 SwRegister_sw_arb_urgent  <= swreg28(9);
 SwRegister_sw_arb_enable  <= swreg28(8);
 SwRegister_sw_arb_time_window_exp  <= swreg28(4 downto 0);
 SwRegister_sw_arb_winer_id  <= swreg29(23 downto 16);
 SwRegister_sw_arb_cur_id  <= swreg29(15 downto 8);
 SwRegister_sw_arb_grp_info  <= swreg29(7 downto 6);
 SwRegister_sw_arb_state  <= swreg29(5 downto 4);
 SwRegister_sw_arb_rst  <= swreg29(3);
 SwRegister_sw_arb_ack  <= swreg29(2);
 SwRegister_sw_arb_fe  <= swreg29(1);
 SwRegister_sw_arb_req  <= swreg29(0);
 SwRegister_sw_arb_satisfaction  <= swreg30(31 downto 0);
