--signal declaration from Document Version v1.5.3
 signal SwRegister_sw_HW_ID : std_logic_vector(15 downto 0);
 signal SwRegister_sw_HW_Version : std_logic_vector(15 downto 0);
 signal SwRegister_sw_HW_BuildDate : std_logic_vector(31 downto 0);
 signal SwRegister_sw_ext_abn_intr_src : std_logic_vector(15 downto 0);
 signal SwRegister_sw_ext_norm_intr_src : std_logic_vector(15 downto 0);
 signal SwRegister_sw_exe_cmdbuf_count : std_logic_vector(31 downto 0);
 signal SwRegister_sw_cmd_exe : std_logic_vector(31 downto 0);
 signal SwRegister_sw_cmd_exe_msb : std_logic_vector(31 downto 0);
 signal SwRegister_sw_axi_TotalARLen : std_logic_vector(31 downto 0);
 signal SwRegister_sw_axi_TotalR : std_logic_vector(31 downto 0);
 signal SwRegister_sw_axi_TotalAR : std_logic_vector(31 downto 0);
 signal SwRegister_sw_axi_TotalRLast : std_logic_vector(31 downto 0);
 signal SwRegister_sw_axi_TotalAWLen : std_logic_vector(31 downto 0);
 signal SwRegister_sw_axi_TotalW : std_logic_vector(31 downto 0);
 signal SwRegister_sw_axi_TotalAW : std_logic_vector(31 downto 0);
 signal SwRegister_sw_axi_TotalWLast : std_logic_vector(31 downto 0);
 signal SwRegister_sw_axi_TotalB : std_logic_vector(31 downto 0);
 signal SwRegister_sw_axi_ARVALID : std_logic;
 signal SwRegister_sw_axi_ARREADY : std_logic;
 signal SwRegister_sw_axi_RVALID : std_logic;
 signal SwRegister_sw_axi_RREADY : std_logic;
 signal SwRegister_sw_axi_AWVALID : std_logic;
 signal SwRegister_sw_axi_AWREADY : std_logic;
 signal SwRegister_sw_axi_WVALID : std_logic;
 signal SwRegister_sw_axi_WREADY : std_logic;
 signal SwRegister_sw_axi_BVALID : std_logic;
 signal SwRegister_sw_axi_BREADY : std_logic;
 signal SwRegister_sw_HW_ApbArbiter : std_logic;
 signal SwRegister_sw_HW_InitMode : std_logic;
 signal SwRegister_sw_core_state : std_logic_vector(4 downto 0);
 signal SwRegister_sw_init_mode : std_logic;
 signal SwRegister_sw_work_state : std_logic_vector(2 downto 0);
 signal SwRegister_sw_arb_check_en : std_logic;
 signal SwRegister_sw_init_enable : std_logic;
 signal SwRegister_sw_axi_clk_gate_disable : std_logic;
 signal SwRegister_sw_master_out_clk_gate_disable : std_logic;
 signal SwRegister_sw_core_clk_gate_disable : std_logic;
 signal SwRegister_sw_abort_mode : std_logic;
 signal SwRegister_sw_reset_core : std_logic;
 signal SwRegister_sw_reset_all : std_logic;
 signal SwRegister_sw_start_trigger : std_logic;
 signal SwRegister_sw_irq_arbrst : std_logic;
 signal SwRegister_sw_irq_jmp : std_logic;
 signal SwRegister_sw_irq_arberr : std_logic;
 signal SwRegister_sw_irq_abort : std_logic;
 signal SwRegister_sw_irq_cmderr : std_logic;
 signal SwRegister_sw_irq_timeout : std_logic;
 signal SwRegister_sw_irq_buserr : std_logic;
 signal SwRegister_sw_irq_endcmd : std_logic;
 signal SwRegister_sw_irq_arbrst_en : std_logic;
 signal SwRegister_sw_irq_jmp_en : std_logic;
 signal SwRegister_sw_irq_arberr_en : std_logic;
 signal SwRegister_sw_irq_abort_en : std_logic;
 signal SwRegister_sw_irq_cmderr_en : std_logic;
 signal SwRegister_sw_irq_timeout_en : std_logic;
 signal SwRegister_sw_irq_buserr_en : std_logic;
 signal SwRegister_sw_irq_endcmd_en : std_logic;
 signal SwRegister_sw_timeout_enable : std_logic;
 signal SwRegister_sw_timeout_cycles : std_logic_vector(30 downto 0);
 signal SwRegister_sw_cmdbuf_exe_addr : std_logic_vector(31 downto 0);
 signal SwRegister_sw_cmdbuf_exe_addr_msb : std_logic_vector(31 downto 0);
 signal SwRegister_sw_cmdbuf_exe_length : std_logic_vector(15 downto 0);
 signal SwRegister_sw_cmd_swap : std_logic_vector(3 downto 0);
 signal SwRegister_sw_data_swap : std_logic_vector(3 downto 0);
 signal SwRegister_sw_max_burst_len : std_logic_vector(7 downto 0);
 signal SwRegister_sw_axi_id_rd : std_logic_vector(7 downto 0);
 signal SwRegister_sw_axi_id_wr : std_logic_vector(7 downto 0);
 signal SwRegister_sw_rdy_cmdbuf_count : std_logic_vector(31 downto 0);
 signal SwRegister_sw_ext_abn_intr_gate : std_logic_vector(15 downto 0);
 signal SwRegister_sw_ext_norm_intr_gate : std_logic_vector(15 downto 0);
 signal SwRegister_sw_cmdbuf_exe_id : std_logic_vector(31 downto 0);
 signal SwRegister_sw_sram_timing_ctrl : std_logic_vector(31 downto 0);
 signal SwRegister_sw_arb_weight : std_logic_vector(4 downto 0);
 signal SwRegister_sw_arb_bw_overflow : std_logic;
 signal SwRegister_sw_arb_urgent : std_logic;
 signal SwRegister_sw_arb_enable : std_logic;
 signal SwRegister_sw_arb_time_window_exp : std_logic_vector(4 downto 0);
 signal SwRegister_sw_arb_winer_id : std_logic_vector(7 downto 0);
 signal SwRegister_sw_arb_cur_id : std_logic_vector(7 downto 0);
 signal SwRegister_sw_arb_grp_info : std_logic_vector(1 downto 0);
 signal SwRegister_sw_arb_state : std_logic_vector(1 downto 0);
 signal SwRegister_sw_arb_rst : std_logic;
 signal SwRegister_sw_arb_ack : std_logic;
 signal SwRegister_sw_arb_fe : std_logic;
 signal SwRegister_sw_arb_req : std_logic;
 signal SwRegister_sw_arb_satisfaction : std_logic_vector(31 downto 0);
